DHCP V2.3.7
R2 4 9 330
R1 4 10 330
R3 4 7 330

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
